** Profile: "SCHEMATIC1-Sweep2"  [ D:\Anselmo\Escritorio\Segundo\FE\Practica4\Apartado1\Ap1-PSpiceFiles\SCHEMATIC1\Sweep2.sim ] 

** Creating circuit file "Sweep2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_Vb 0 1 0.001 
.STEP LIN V_Vce 0 20 5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
