** Profile: "SCHEMATIC1-Practica6_3"  [ C:\Users\juanc\Desktop\Teleco\Segundo\FE\Practica6\Practica6_3-PSpiceFiles\SCHEMATIC1\Practica6_3.sim ] 

** Creating circuit file "Practica6_3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../practica6_3-pspicefiles/practica6_3.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 5us 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
