** Profile: "SCHEMATIC1-sweep"  [ D:\Anselmo\Escritorio\Segundo\FE\Practica4\Apartado1\Ap1-PSpiceFiles\SCHEMATIC1\sweep.sim ] 

** Creating circuit file "sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_Vce 0 10 0.01 
.STEP LIN I_Ib 0 100uA 10uA 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
